module trajectory_mif_writer(
	trajectory_memloc,
	trajectory_memloc_enable,
	rd_add(character_address),
	rd_clk(character_clock),
	rd_out(character_out)
);

endmodule
