module ascii_to_number (ascii, number);

	input[47:0] ascii;
	output[31:0] number;
	
	reg[31:0] ones, tens, hundreds, thousands, tenth, hundth;
	always @(ascii)
	begin
		ones <= 
	end
		
endmodule
